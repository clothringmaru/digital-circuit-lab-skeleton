`ifndef __ALUFUNC_VH__
`define __ALUFUNC_VH__

`define ALU_ADD     3'b000
`define ALU_SUB     3'b001
`define ALU_AND     3'b010
`define ALU_OR      3'b011
`define ALU_MOVI        3'b100      
`endif
